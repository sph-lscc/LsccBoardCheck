/* synthesis translate_off*/
`define SIM
/* synthesis translate_on*/
`ifndef SIM
`define SYNTH
`endif

`timescale 1 ns / 1 ps
